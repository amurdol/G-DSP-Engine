// ============================================================================
// G-DSP Engine — System Top-Level
// ============================================================================
// Author : G-DSP Team
// Project: TFG — 16-QAM Baseband Processor on Gowin GW1NR-9
// License: MIT
// ============================================================================
//
// Top-level integration for Sipeed Tang Nano 9K:
//
//   ┌─────────────────────────────────────────────────────────────────────┐
//   │  clk_27m (27 MHz)                                                   │
//   │      │                                                              │
//   │      ▼                                                              │
//   │  ┌───────┐   clk_dsp (27 MHz)                                       │
//   │  │ GW_PLL├──────────────────┐                                       │
//   │  │       │   clk_pixel (25.2 MHz, VGA 480p)                         │
//   │  │       ├────────────────┐ │                                       │
//   │  │       │   clk_serial (126 MHz)                                   │
//   │  │       ├──────────────┐ │ │                                       │
//   │  └───────┘              │ │ │                                       │
//   │                         │ │ │                                       │
//   │  ┌─────────┐  ┌─────────┴─┴─┴───────────────────────────────────┐   │
//   │  │         │  │ clk_dsp domain                                  │   │
//   │  │  Button │  │  tx_top → channel_top → rx_top                  │   │
//   │  │   S1    │──│    (PRBS→QAM→RRC→AWGN→RRC→Gardner→Costas)      │   │
//   │  │         │  │                                    ↓            │   │
//   │  └─────────┘  │                             demod_I/Q/valid     │   │
//   │               └──────────────────────────────────────┬──────────┘   │
//   │                                                      │              │
//   │               ┌──────────────────────────────────────┼──────────┐   │
//   │               │ clk_pixel domain                     ↓          │   │
//   │               │  constellation_renderer → hdmi_tx → TMDS       │   │
//   │               │  (640×480 @ 60 Hz VGA)                          │   │
//   │               └────────────────────────────────────────────────┘   │
//   └─────────────────────────────────────────────────────────────────────┘
//
// Button S1 cycles diagnostic display mode:
//   Mode 0: QAM mapper output (raw symbols → expect 16 clean points)
//   Mode 1: TX RRC output (post pulse-shaping → ISI visible)
//   Mode 2: Channel output (TX + noise)
//   Mode 3: Full RX chain (through Costas loop demod)
// LEDs[2:3] display current mode, LED[1]=lock, LED[4]=PLL, LED[5]=heartbeat
// ============================================================================

module gdsp_top
    import gdsp_pkg::*;
(
    input  logic        clk_27m,        // 27 MHz board oscillator
    input  logic        rst_n,          // Active-low reset (button S2)
    input  logic        btn_user,       // User button S1 (noise control)
    output logic [5:0]  led,            // Onboard LEDs (active-low)

    // --- HDMI TMDS output (differential via ELVDS_OBUF) ---
    output logic        tmds_clk_p,
    output logic        tmds_clk_n,
    output logic [2:0]  tmds_data_p,
    output logic [2:0]  tmds_data_n
);

    // ========================================================================
    // Clock Generation for VGA 480p HDMI
    //
    // Architecture:
    //   clk_27m (27 MHz)
    //       │
    //       ├──────────────────────────────► clk_dsp (27 MHz, direct)
    //       │
    //       ▼
    //   ┌─────────┐   clk_serial (126 MHz)
    //   │Gowin_rPLL├────────────────────────► to HDMI serialiser (5× pixel)
    //   │         │         │
    //   └─────────┘         ▼
    //               ┌────────────┐
    //               │Gowin_CLKDIV│  ÷5
    //               │            ├──────────► clk_pixel (25.2 MHz, VGA 480p)
    //               └────────────┘
    //
    // PLL Config: VCO = 27×14/3 = 126 MHz, CLKOUT = 126 MHz
    //             (IDIV=2 [÷3], FBDIV=13 [×14], ODIV=4 [÷4])
    // ========================================================================
    logic clk_dsp;
    logic clk_pixel;
    logic clk_serial;
    logic pll_lock;

    // DSP clock = input clock directly (27 MHz)
    assign clk_dsp = clk_27m;

    // rPLL: 27 MHz → 126 MHz (clk_serial for VGA 480p HDMI TMDS)
    // VCO = 27×14/3 = 126 MHz, ODIV divides by 4
    // Hardware: IDIV=2 (÷3), FBDIV=13 (×14), ODIV=4 (÷4)
    Gowin_rPLL u_pll (
        .clkin  (clk_27m),
        .clkout (clk_serial),    // 126 MHz (5× pixel clock)
        .lock   (pll_lock)
    );

    // CLKDIV: 126 MHz ÷ 5 → 25.2 MHz (VGA 480p pixel clock)
    Gowin_CLKDIV u_clkdiv (
        .hclkin (clk_serial),
        .resetn (pll_lock),      // Hold in reset until PLL locks
        .clkout (clk_pixel)      // 25.2 MHz
    );

    // Combined reset: external button AND PLL lock
    wire sys_rst_n = rst_n && pll_lock;

    // ========================================================================
    // Button Debouncer + Noise Level Cycler (S1)
    //
    // Debounce: ~20ms at 27 MHz ≈ 540,000 cycles → use 19-bit counter
    // Noise levels: 0 → 20 → 50 → 100 (cycle on press)
    // ========================================================================
    logic [18:0] debounce_cnt;
    logic        btn_sync0, btn_sync1, btn_stable, btn_prev;
    logic [1:0]  noise_sel;
    logic [NOISE_MAG_WIDTH-1:0] noise_magnitude;

    // Synchroniser
    always_ff @(posedge clk_dsp or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            btn_sync0 <= 1'b1;  // Default high (button released)
            btn_sync1 <= 1'b1;
        end else begin
            btn_sync0 <= btn_user;
            btn_sync1 <= btn_sync0;
        end
    end

    // Debounce counter
    always_ff @(posedge clk_dsp or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            debounce_cnt <= '0;
            btn_stable   <= 1'b1;
        end else begin
            if (btn_sync1 != btn_stable) begin
                if (debounce_cnt == 19'h7FFFF)
                    btn_stable <= btn_sync1;
                else
                    debounce_cnt <= debounce_cnt + 1'b1;
            end else begin
                debounce_cnt <= '0;
            end
        end
    end

    // Edge detect for button press (falling edge = button pressed)
    always_ff @(posedge clk_dsp or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            btn_prev  <= 1'b1;
            noise_sel <= 2'b00;
        end else begin
            btn_prev <= btn_stable;
            if (btn_prev && !btn_stable)  // Falling edge
                noise_sel <= noise_sel + 1'b1;
        end
    end

    // Diagnostic mode: noise fixed to 0 for clean bypass testing
    assign noise_magnitude = 8'd0;

    // ========================================================================
    // TX Subsystem
    // ========================================================================
    sample_t tx_I, tx_Q;
    logic    tx_valid;
    logic    sym_tick;
    sample_t map_I, map_Q;
    logic    map_valid;

    tx_top u_tx (
        .clk       (clk_dsp),
        .rst_n     (sys_rst_n),
        .en        (1'b1),
        .tx_I      (tx_I),
        .tx_Q      (tx_Q),
        .tx_valid  (tx_valid),
        .sym_tick  (sym_tick),
        .map_I     (map_I),
        .map_Q     (map_Q),
        .map_valid (map_valid)
    );

    // ========================================================================
    // AWGN Channel
    // ========================================================================
    sample_t ch_I, ch_Q;
    logic    ch_valid;

    channel_top u_channel (
        .clk             (clk_dsp),
        .rst_n           (sys_rst_n),
        .en              (1'b1),
        .tx_I            (tx_I),
        .tx_Q            (tx_Q),
        .tx_valid        (tx_valid),
        .noise_magnitude (noise_magnitude),
        .rx_I            (ch_I),
        .rx_Q            (ch_Q),
        .rx_valid        (ch_valid)
    );

    // ========================================================================
    // RX Subsystem
    // ========================================================================
    sample_t demod_I, demod_Q;
    logic    demod_valid;
    logic    demod_lock;

    rx_top u_rx (
        .clk         (clk_dsp),
        .rst_n       (sys_rst_n),
        .rx_I        (ch_I),
        .rx_Q        (ch_Q),
        .rx_valid    (ch_valid),
        .demod_I     (demod_I),
        .demod_Q     (demod_Q),
        .demod_valid (demod_valid),
        .demod_lock  (demod_lock)
    );

    // ========================================================================
    // Diagnostic Display Mux
    //
    // Button S1 (noise_sel) selects which signal feeds the renderer:
    //   0 = QAM mapper symbols (raw, pre-RRC)   → expect 16 clean dots
    //   1 = TX output (post-RRC pulse shaping)   → ISI visible
    //   2 = Channel output (TX + noise)          → noise = 0 for diag
    //   3 = RX demod output (after Costas loop)  → normal operation
    // ========================================================================
    sample_t disp_I, disp_Q;
    logic    disp_valid;

    always_comb begin
        case (noise_sel)
            2'b00: begin
                disp_I     = map_I;
                disp_Q     = map_Q;
                disp_valid = map_valid;
            end
            2'b01: begin
                disp_I     = tx_I;
                disp_Q     = tx_Q;
                disp_valid = tx_valid & sym_tick;  // Gate to symbol rate
            end
            2'b10: begin
                disp_I     = ch_I;
                disp_Q     = ch_Q;
                disp_valid = ch_valid & sym_tick;  // Gate to symbol rate
            end
            2'b11: begin
                disp_I     = demod_I;
                disp_Q     = demod_Q;
                disp_valid = demod_valid;
            end
            default: begin
                disp_I     = demod_I;
                disp_Q     = demod_Q;
                disp_valid = demod_valid;
            end
        endcase
    end

    // ========================================================================
    // Constellation Renderer (clk_pixel domain)
    //
    // sym_valid from DSP domain needs CDC — the renderer handles this
    // internally with a 2-FF synchroniser.
    // ========================================================================
    logic [23:0] rgb_pixel;
    logic        video_hsync, video_vsync, video_de;

    constellation_renderer u_renderer (
        .clk_pixel  (clk_pixel),
        .rst_n      (sys_rst_n),
        .sym_I      (disp_I),
        .sym_Q      (disp_Q),
        .sym_valid  (disp_valid),
        .rgb_pixel  (rgb_pixel),
        .hsync      (video_hsync),
        .vsync      (video_vsync),
        .de         (video_de)
    );

    // ========================================================================
    // HDMI Transmitter (TMDS encoding + serialisation)
    // ========================================================================
    hdmi_tx u_hdmi (
        .clk_pixel  (clk_pixel),
        .clk_serial (clk_serial),
        .rst_n      (sys_rst_n),
        .rgb        (rgb_pixel),
        .hsync      (video_hsync),
        .vsync      (video_vsync),
        .de         (video_de),
        .tmds_clk_p (tmds_clk_p),
        .tmds_clk_n (tmds_clk_n),
        .tmds_d_p   (tmds_data_p),
        .tmds_d_n   (tmds_data_n)
    );

    // ========================================================================
    // LED Indicators (active-low) - NO dependen de PLL lock para debug
    //
    // LED[0]: Heartbeat (~0.8 Hz blink) - usa rst_n directo
    // LED[1]: PLL lock status (lit = locked)
    // LED[2]: Costas lock indicator (lit = locked)
    // LED[3]: sys_rst_n status (lit = system running)
    // LED[4]: Noise level bit 0
    // LED[5]: Noise level bit 1
    // ========================================================================
    logic [24:0] heartbeat_cnt;

    // Heartbeat usa rst_n directo, NO sys_rst_n
    always_ff @(posedge clk_dsp or negedge rst_n) begin
        if (!rst_n)
            heartbeat_cnt <= '0;
        else
            heartbeat_cnt <= heartbeat_cnt + 1'b1;
    end

    // LED mapping (active-low, per design spec):
    // LED[0]: reset status
    // LED[1]: demodulator lock (Costas loop phase lock)
    // LED[2-3]: diagnostic display mode (00=mapper, 01=TX, 10=ch, 11=demod)
    // LED[4]: PLL lock
    // LED[5]: heartbeat
    assign led[0] = ~sys_rst_n;           // Reset indicator (active-low)
    assign led[1] = ~demod_lock;          // Demod lock status
    assign led[2] = ~noise_sel[0];        // Diag mode bit 0
    assign led[3] = ~noise_sel[1];        // Diag mode bit 1
    assign led[4] = ~pll_lock;            // PLL lock diagnostic
    assign led[5] = ~heartbeat_cnt[24];   // Heartbeat (must always blink)

endmodule : gdsp_top

// ============================================================================
// Gowin IP Simulation Stubs
//
// These modules are ONLY for Icarus Verilog simulation.
// For Gowin synthesis, the actual IPs in src/gowin_rpll/ and src/gowin_clkdiv/
// are used instead.
// ============================================================================
`ifdef SIMULATION

module Gowin_rPLL (
    input  logic clkin,
    output logic clkout,
    output logic lock
);
    // Simulation model: generate 126 MHz from 27 MHz input
    assign lock = 1'b1;

    // Generate clk_serial (126 MHz) — period 7.936 ns
    logic clk_ser_sim = 0;
    always #3.968 clk_ser_sim = ~clk_ser_sim;
    assign clkout = clk_ser_sim;
endmodule : Gowin_rPLL

module Gowin_CLKDIV (
    input  logic hclkin,
    input  logic resetn,
    output logic clkout
);
    // Simulation model: divide input by 5
    // 126 MHz / 5 = 25.2 MHz — period 39.68 ns
    logic clk_pix_sim = 0;
    always #19.84 clk_pix_sim = ~clk_pix_sim;
    assign clkout = resetn ? clk_pix_sim : 1'b0;
endmodule : Gowin_CLKDIV

// OSER10: 10:1 Serialiser (simulation stub — just outputs LSB)
module OSER10 (
    input  logic D0, D1, D2, D3, D4, D5, D6, D7, D8, D9,
    input  logic PCLK,
    input  logic FCLK,
    input  logic RESET,
    output logic Q
);
    // Simulation: just output D0 (LSB) for basic functionality check
    assign Q = D0;
endmodule

// ELVDS_OBUF: LVDS output buffer (simulation stub — passthrough)
module ELVDS_OBUF (
    input  logic I,
    output logic O,
    output logic OB
);
    assign O  = I;
    assign OB = ~I;
endmodule

`endif // SIMULATION
