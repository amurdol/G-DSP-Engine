// Placeholder — RRC FIR pulse-shaping / matched filter
// To be implemented in Phase 1
