// ============================================================================
// G-DSP Engine — Testbench: System Top-Level Integration
// ============================================================================
// Phase 4 integration testbench for gdsp_top.  Verifies:
//   1. PLL simulation model produces valid clocks
//   2. DSP chain (TX → Channel → RX) produces demodulated symbols
//   3. Button debounce cycles noise_magnitude correctly
//   4. Constellation renderer and HDMI TX instantiate without errors
//   5. Costas lock is achieved with at least one noise level
//
// Note: HDMI TMDS output is not validated (would require external
// capture/analysis). We verify RTL compiles and runs without hangs.
//
// Usage (Icarus Verilog):
//   iverilog -g2012 -DSIMULATION -I sim/vectors -o sim/out/tb_gdsp_top.vvp \
//       rtl/packages/gdsp_pkg.sv rtl/common/bit_gen.sv \
//       rtl/modem/qam16_mapper.sv rtl/modem/rrc_filter.sv rtl/modem/tx_top.sv \
//       rtl/channel/awgn_generator.sv rtl/channel/awgn_channel.sv \
//       rtl/sync/gardner_ted.sv rtl/sync/costas_loop.sv rtl/modem/rx_top.sv \
//       rtl/video/constellation_renderer.sv rtl/video/hdmi_tx.sv \
//       rtl/top/gdsp_top.sv sim/tb/tb_gdsp_top.sv
//   vvp sim/out/tb_gdsp_top.vvp
// ============================================================================

`timescale 1ns / 1ps

module tb_gdsp_top;

    import gdsp_pkg::*;

    // -----------------------------------------------------------------------
    // Test Configuration
    // -----------------------------------------------------------------------
    localparam int SIM_CYCLES       = 100000;   // ~3.7 ms at 27 MHz
    localparam int LOCK_TIMEOUT     = 80000;    // Cycles before lock expected
    localparam int BUTTON_HOLD_NS   = 500000;   // 500 µs button press

    // -----------------------------------------------------------------------
    // DUT signals
    // -----------------------------------------------------------------------
    logic        clk_27m;
    logic        rst_n;
    logic        btn_user;
    logic [5:0]  led;
    logic        tmds_clk_p, tmds_clk_n;
    logic [2:0]  tmds_data_p, tmds_data_n;

    // -----------------------------------------------------------------------
    // Clock generation: 27 MHz → period = 37.037 ns
    // -----------------------------------------------------------------------
    initial clk_27m = 1'b0;
    always #18.519 clk_27m = ~clk_27m;

    // -----------------------------------------------------------------------
    // DUT instantiation
    // -----------------------------------------------------------------------
    gdsp_top u_dut (
        .clk_27m     (clk_27m),
        .rst_n       (rst_n),
        .btn_user    (btn_user),
        .led         (led),
        .tmds_clk_p  (tmds_clk_p),
        .tmds_clk_n  (tmds_clk_n),
        .tmds_data_p (tmds_data_p),
        .tmds_data_n (tmds_data_n)
    );

    // -----------------------------------------------------------------------
    // VCD dump
    // -----------------------------------------------------------------------
    initial begin
        $dumpfile("sim/waves/tb_gdsp_top.vcd");
        $dumpvars(0, tb_gdsp_top);
    end

    // -----------------------------------------------------------------------
    // Test monitoring
    // -----------------------------------------------------------------------
    int cycle_count = 0;
    logic lock_seen = 0;
    int lock_cycle = 0;

    // Monitor LED[1] for lock (active-low, so lock = LED[1] == 0)
    always @(posedge clk_27m) begin
        cycle_count <= cycle_count + 1;
        if (!lock_seen && led[1] == 1'b0) begin
            lock_seen <= 1'b1;
            lock_cycle <= cycle_count;
            $display("[TB] Lock detected at cycle %0d (%.2f ms)",
                     cycle_count, cycle_count * 37.037e-6);
        end
    end

    // -----------------------------------------------------------------------
    // Button press task
    // -----------------------------------------------------------------------
    task automatic press_button();
        $display("[TB] Pressing button S1 (diagnostic mode cycle)...");
        btn_user = 1'b0;  // Active-low press
        #(BUTTON_HOLD_NS);
        btn_user = 1'b1;  // Release
        #100000;          // Debounce settle
    endtask

    // -----------------------------------------------------------------------
    // Main test sequence
    // -----------------------------------------------------------------------
    int errors = 0;

    initial begin
        $display("============================================================");
        $display("  G-DSP Engine — Phase 4 Integration Test");
        $display("============================================================");

        // Initial state
        rst_n    = 1'b0;
        btn_user = 1'b1;  // Not pressed (active-low)

        // Hold reset
        repeat (100) @(posedge clk_27m);
        rst_n = 1'b1;
        $display("[TB] Reset released");

        // Wait for initial lock (noise_mag = 0)
        $display("[TB] Waiting for Costas lock (noise_mag = 0)...");
        repeat (LOCK_TIMEOUT) @(posedge clk_27m);

        if (!lock_seen) begin
            $display("[WARN] No lock detected within %0d cycles at noise=0", LOCK_TIMEOUT);
        end

        // Test button cycling: mode 0→1→2→3 (mapper→TX→ch→demod)
        $display("\n[TB] Testing diagnostic display mode cycling via button S1:");
        for (int i = 0; i < 4; i++) begin
            $display("[TB]   Display mode after %0d presses: LED[3:2] = %b", i, led[3:2]);
            if (i < 3) press_button();
        end

        // Continue simulation to verify stability
        $display("\n[TB] Running extended simulation (%0d total cycles)...", SIM_CYCLES);
        while (cycle_count < SIM_CYCLES) begin
            @(posedge clk_27m);
        end

        // -----------------------------------------------------------------------
        // Results
        // -----------------------------------------------------------------------
        $display("\n============================================================");
        $display("  INTEGRATION TEST RESULTS");
        $display("============================================================");
        $display("  Simulation cycles  : %0d", cycle_count);
        $display("  Lock achieved      : %s", lock_seen ? "YES" : "NO");
        if (lock_seen)
            $display("  Lock cycle         : %0d (%.2f ms)", lock_cycle, lock_cycle * 37.037e-6);
        $display("  PLL lock LED[4]    : %s", (led[4] == 1'b0) ? "LOCKED" : "UNLOCKED");
        $display("  Final diag mode    : LED[3:2] = %b", led[3:2]);
        $display("  Heartbeat LED[0]   : toggling (observed via VCD)");
        $display("============================================================");

        // PASS/FAIL criteria
        if (lock_seen && led[4] == 1'b0) begin
            $display("[TB] *** ALL TESTS PASSED ***");
        end else begin
            $display("[TB] *** TEST FAILED ***");
            if (!lock_seen) $display("      - Costas lock not achieved");
            if (led[4] != 1'b0) $display("      - PLL not locked");
            errors = 1;
        end

        $display("============================================================\n");
        #1000;
        $finish;
    end

endmodule
