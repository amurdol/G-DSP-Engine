// ============================================================================
// G-DSP Engine — Root-Raised Cosine (RRC) FIR Filter
// ============================================================================
// 33-tap symmetric FIR filter implementing pulse shaping (Tx) or matched
// filtering (Rx) for the 16-QAM modem.
//
// Architecture: **Transposed-Form FIR**
//
//   Why transposed form?
//   1. Each tap = one multiplier + one adder + one register.  The register
//      sits at the output of each stage, which maps directly onto the
//      Gowin pREG+MULT9 primitive (DSP slice post-multiply register).
//   2. The critical path is a single multiply + add, regardless of the
//      number of taps.  This is the shortest achievable for FIR.
//   3. No long accumulator chain — the additions are distributed.
//
//   Why NOT folded/time-multiplexed?
//   At 27 MHz system clock with SPS=4, the sample rate is 27 MHz.
//   A folded architecture for 33 taps would need 33 multiply cycles per
//   sample → 33 x 27 MHz = 891 MHz internal clock.  Impossible on GW1NR-9.
//   The transposed form processes one sample per clock at 27 MHz.
//
//   DSP budget: 33 taps × 2 (I+Q) = 66 multipliers.  The GW1NR-9 has 20
//   MULT9 slices (= 10 MULT18).  Since 12×12 requires MULT18 mode, we
//   would need 33 MULT18 per channel → not enough for fully parallel.
//
//   **Symmetry exploitation**: The RRC filter has linear-phase symmetry
//   (h[n] = h[N-1-n]).  We fold symmetric taps: add x[n]+x[N-1-n] BEFORE
//   multiplying → only ceil(33/2) = 17 multipliers per channel.
//   Two channels (I+Q) = 34 multipliers @ MULT18 → still 34 > 10.
//
//   **Practical compromise**: We use transposed form with fabric multipliers.
//   The Gowin synthesiser will map as many multiplies as possible into the
//   available MULT9/MULT18 slices and implement the rest in LUT-based
//   multipliers.  At 12×12 bits and 27 MHz, LUT-based multipliers will
//   easily meet timing.  Resource estimate: ~33 × ~144 LUT4 ≈ 4,752 LUTs
//   per channel.  With both I and Q sharing the same coefficient set, total
//   ≈ 9,504 LUTs — tight for 8,640 LUTs.
//
//   **FINAL DECISION — Folded with dual-clock trick is unrealistic.**
//   **We use transposed form for a SINGLE channel; tx_top instantiates
//   TWO rrc_filter instances (I and Q).  DSP slices will be shared by
//   Gowin's resource-sharing pass.  If resource pressure is too high we
//   will time-multiplex I/Q in Phase 4 (integration).**
//
// Coefficient loading:
//   Coefficients are loaded from an `include` file generated by the
//   Python Golden Model (sim/vectors/rrc_coeffs.v).
//
// Data flow:
//   din (Q1.11) --[×coeff]-- → product (Q2.22, 24-bit) → truncate → dout
//
// Latency: NUM_TAPS clock cycles (fully pipelined, 1 output per clock)
// ============================================================================

module rrc_filter
    import gdsp_pkg::*;
(
    input  logic     clk,
    input  logic     rst_n,
    input  sample_t  din,       // Input sample  (Q1.11, 12-bit signed)
    input  logic     din_valid, // Input valid strobe
    output sample_t  dout,      // Filtered output (Q1.11, 12-bit signed)
    output logic     dout_valid // Output valid strobe
);

    // -----------------------------------------------------------------------
    // Coefficient ROM — loaded from auto-generated include file
    // -----------------------------------------------------------------------
    `include "../../sim/vectors/rrc_coeffs.v"
    // Provides: localparam signed [11:0] RRC_COEFFS [0:32]

    // -----------------------------------------------------------------------
    // Transposed FIR pipeline registers
    //
    //  Stage N-1:  product[N-1] = din * coeff[N-1]
    //  Stage k  :  pipe[k]      = din * coeff[k] + pipe[k+1]
    //  Output   :  dout         = pipe[0] (truncated to 12 bits)
    //
    //  We use ACCUM_WIDTH (30 bits) for the pipeline registers to prevent
    //  any overflow during accumulation.  The products are 24 bits but we
    //  sign-extend to 30 bits before adding.
    // -----------------------------------------------------------------------

    // Product wires (combinational multiply)
    logic signed [PRODUCT_WIDTH-1:0] product [0:NUM_TAPS-1];

    // Transposed pipeline registers
    logic signed [ACCUM_WIDTH-1:0] pipe_r [0:NUM_TAPS-1];

    // Valid delay line (match pipeline latency = 1 cycle for transposed)
    logic valid_d1;

    // -----------------------------------------------------------------------
    // Combinational: multiply input by each coefficient
    //   Structured as:  product = din * coeff
    //   The synthesiser will infer MULT18 or LUT multipliers.
    // -----------------------------------------------------------------------
    always_comb begin
        for (int i = 0; i < NUM_TAPS; i++) begin
            product[i] = din * RRC_COEFFS[i];
        end
    end

    // -----------------------------------------------------------------------
    // Sequential: transposed-form pipeline
    //   pipe[N-1] = product[N-1]                    (last stage, no add)
    //   pipe[k]   = product[k] + pipe[k+1]_prev     (k = N-2 downto 0)
    //   Output is pipe[0] after truncation.
    // -----------------------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int i = 0; i < NUM_TAPS; i++) begin
                pipe_r[i] <= '0;
            end
            valid_d1 <= 1'b0;
        end else begin
            valid_d1 <= din_valid;
            if (din_valid) begin
                // Last stage: just the product (sign-extended to ACCUM_WIDTH)
                pipe_r[NUM_TAPS-1] <= ACCUM_WIDTH'(product[NUM_TAPS-1]);

                // Remaining stages: product + previous pipe value from next stage
                for (int i = 0; i < NUM_TAPS-1; i++) begin
                    pipe_r[i] <= ACCUM_WIDTH'(product[i]) + pipe_r[i+1];
                end
            end
        end
    end

    // -----------------------------------------------------------------------
    // Output truncation with convergent rounding
    //
    //   pipe_r[0] is in Q format:
    //     Input  = Q1.11 (12-bit), Coeff = Q1.11 (12-bit)
    //     Product = Q2.22 (24-bit), sign-extended to 30 bits
    //     After accumulation: still Q2.22 in 30 bits (symmetric filter,
    //       sum of |coeff| < 1, so no integer overflow)
    //
    //   To truncate back to Q1.11 (12-bit output):
    //     - Discard the top guard bits (keep from bit 22 downward)
    //     - Keep 12 bits: [22:11] gives Q1.11
    //     - Bits [10:0] are the truncated fractional bits
    //
    //   Convergent (banker's) rounding:
    //     round_bit  = pipe_r[0][10]         (MSB of truncated portion)
    //     sticky_bits = |pipe_r[0][9:0]      (OR of remaining)
    //     round_up = round_bit & (sticky_bits | pipe_r[0][11])
    //                                         (round to even)
    // -----------------------------------------------------------------------
    logic signed [ACCUM_WIDTH-1:0] acc_val;
    logic round_bit, sticky, lsb_result;
    logic round_up;
    sample_t dout_trunc;

    assign acc_val    = pipe_r[0];
    assign round_bit  = acc_val[FRAC_BITS-1];              // bit [10]
    assign sticky     = |acc_val[FRAC_BITS-2:0];           // bits [9:0]
    assign lsb_result = acc_val[FRAC_BITS];                // bit [11]
    assign round_up   = round_bit & (sticky | lsb_result); // convergent

    // Truncate: take bits [22:11] and add rounding
    assign dout_trunc = acc_val[FRAC_BITS + DATA_WIDTH - 1 : FRAC_BITS]
                        + {{(DATA_WIDTH-1){1'b0}}, round_up};

    // -----------------------------------------------------------------------
    // Saturation check (safety — should never trigger with properly
    // normalised coefficients, but protects against unexpected overflow)
    // -----------------------------------------------------------------------
    localparam sample_t SAT_POS =  (1 <<< (DATA_WIDTH-1)) - 1;  // +2047
    localparam sample_t SAT_NEG = -(1 <<< (DATA_WIDTH-1));       // -2048

    sample_t dout_sat;

    always_comb begin
        // Check if the upper bits (above bit 22) carry meaningful magnitude
        // If acc_val[ACCUM_WIDTH-1:FRAC_BITS+DATA_WIDTH-1] are not all the
        // same (sign extension), then we have overflow.
        if (acc_val[ACCUM_WIDTH-1] == 1'b0 &&
            |acc_val[ACCUM_WIDTH-1 : FRAC_BITS+DATA_WIDTH] != 1'b0) begin
            dout_sat = SAT_POS;   // Positive overflow
        end else if (acc_val[ACCUM_WIDTH-1] == 1'b1 &&
                     &acc_val[ACCUM_WIDTH-1 : FRAC_BITS+DATA_WIDTH] != 1'b1) begin
            dout_sat = SAT_NEG;   // Negative overflow
        end else begin
            dout_sat = dout_trunc;
        end
    end

    assign dout       = dout_sat;
    assign dout_valid = valid_d1;

endmodule : rrc_filter
